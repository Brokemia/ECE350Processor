module UART_tb();
    reg clk = 1'b0;
    reg serialIn = 1'b1;
    wire serialOut;
    reg setAddr = 1'b0;
    reg [11:0] startAddr = 12'b0;
    wire err;
    wire [11:0] writeAddr;
    wire [31:0] writeData;
    wire writeEnable;
    UART uut(clk, serialIn, serialOut, setAddr, startAddr, err, writeAddr, writeData, writeEnable);
    initial begin
        $dumpfile("uart.vcd");
        $dumpvars(0, UART_tb);
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        serialIn <= 1'b1;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        clk = 1'b0;
        #10;
        clk = 1'b1;
        #10;
        $finish;
    end
endmodule